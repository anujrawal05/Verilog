module gain_stage(
    input wire clk,
    input wire signed [15:0] input_signal,
    output reg signed [15:0] amplified_output
);

    parameter GAIN = 100;  // Open loop gain
    wire signed [31:0] temp_output;
    
    assign temp_output = input_signal * GAIN;
    
    always @(posedge clk) begin
        // Limit to 16-bit range
        if (temp_output > 32767)
            amplified_output <= 16'd32767;
        else if (temp_output < -32768)
            amplified_output <= -16'd32768;
        else
            amplified_output <= temp_output[15:0];
    end

endmodule 